module tb_dso_board();

endmodule
